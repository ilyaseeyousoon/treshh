module mlt_x400 (input clk, input rst, input[9:0] int_data[7:0], input[6:0] frac_data[7:0], input start, 
					  output[19:0] out_16, output out_dval);

logic[6:0] frac_delay[7:0];
logic[15:0] mult_out[7:0];
logic[16:0] sum_st_1[7:0];
logic[17:0] sum_st_2[3:0];
logic[18:0] sum_st_3[1:0];
logic[19:0] sum_st_4;
logic[4:0] lr_ena;
					  
genvar g;
generate
	for(g = 0; g < 8; g++) begin : gen_mult
		mult_x50 mlt_inst (~rst, start, clk, int_data[g], mult_out[g]);
	end
endgenerate

assign out_dval = lr_ena[4];
assign out_16 = sum_st_4;

integer i;

always_ff @ (posedge clk or negedge rst)
	begin
		if(!rst)
			begin
				lr_ena <= 0;
			end
		else
			begin
				lr_ena <= {lr_ena[3:0], start};
				for(i = 0; i < 8; i++)
					begin
						frac_delay[i] <= (start) ? frac_data[i] : 0;
						sum_st_1[i] <= (lr_ena[0]) ? (mult_out[i] + frac_delay[i]) : 0;
					end
					
				for(i = 0; i < 4; i++)
					sum_st_2[i] <= (lr_ena[1]) ? (sum_st_1[i*2] + sum_st_1[i*2+1]) : 0;
					
				for(i = 0; i < 2; i++)
					sum_st_3[i] <= (lr_ena[2]) ? (sum_st_2[i*2] + sum_st_2[i*2+1]) : 0;
					
				//sum_st_4 <= (lr_ena[3]) ? (sum_st_3[0] + sum_st_3[1]) : 0;
				sum_st_4 <= (sum_st_3[0] + sum_st_3[1]);
				
			end
	end
	
endmodule
	
